module Lab1(input logic a, b, output logic y);
assign y = a & b; // a 2-input digital AND gate
endmodule